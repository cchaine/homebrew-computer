----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:31:09 04/13/2021 
-- Design Name: 
-- Module Name:    counter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity counter is
    Generic (Size : integer := 16);
    Port ( CLK : in  STD_LOGIC;
           RST : in STD_LOGIC;
           OE : in STD_LOGIC;
           CEN : in  STD_LOGIC;
           DIR : in  STD_LOGIC;
           LOAD : in  STD_LOGIC;
           B_Addr : inout  STD_LOGIC_VECTOR (Size-1 downto 0));
end counter;

architecture Behavioral of counter is
   signal value : STD_LOGIC_VECTOR (Size-1 downto 0) := (others => '0');
begin
   B_Addr <= value when OE = '1' else (others => 'Z');
   
   process(RST, CLK)
   begin
      if rising_edge(CLK) then
        -- Counting feature
        if CEN = '1' then
          if DIR = '0' then
            value <= value - 1;
          else
            value <= value + 1;
          end if;
        end if;
        -- Parallel loading feature
        if LOAD = '1' and OE /= '1' then
          value <= B_Addr;
        end if;
      end if;
      -- Asynchronous reset feature
      if rising_edge(RST) then
         value <= (others => '0');
      end if;
   end process;

end Behavioral;

